`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   12:05:11 07/14/2011
// Design Name:   cs_component
// Module Name:   C:/Users/epoxytheory/Documents/CarrierSense/cs_component_tb.v
// Project Name:  CarrierSense
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: cs_component
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module cs_component_tb;

	// Inputs
	reg clk;
	reg rst;
	reg [15:0] real_value;
	reg [15:0] img_value	;
	reg [31:0] count;
	reg run;
	reg done;
	
	wire strobe;
	wire attempt_sample_write;
	wire present;
	wire [15:0] present_nextcount;

	// Instantiate the Unit Under Test (UUT)
	cs_component uut (
		.clk(clk), 
		.rst(rst), 
		.real_value(real_value), 
		.img_value(img_value), 
		.present_next(present),
		.strobe(strobe),
		.run(run),
		.present_nextcount(present_nextcount)
	);
cic_strober cic_strober(.clock(clk),.reset(rst),.enable(1'b1),.rate(320),
			   .strobe_fast(1),.strobe_slow(strobe) ); //strober gives pulse at every 320 clock cycles

	initial begin
		// Initialize Inputs
		clk = 0;
		rst = 0;
		real_value = 0;
		img_value = 0;
		count = 0;
		
		@(posedge clk)
		rst = 1;
		@(posedge clk)
		rst = 0;
		//Wait 100 ns for global reset to finish
		//#100;  
		//Add stimulus here

	end
	
	always begin
	#7.8125 clk = ~clk; //64 MHz clock signal generated by on-board fpga clock
	end

always @(posedge strobe) begin //wait for the strobe to go high
	real_value = $random()%32768; //produce I and Q values for the carrier sense module
	img_value = $random()%32768; 
end

always @ ( posedge strobe) count = count + 1;

      
endmodule

